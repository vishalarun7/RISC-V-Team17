module hazard_unit #(
    
)